module renderer


